library verilog;
use verilog.vl_types.all;
entity memory_tex_vlg_vec_tst is
end memory_tex_vlg_vec_tst;
